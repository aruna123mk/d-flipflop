
`include "dff_seqitm.sv"   // Defines sequence item class
`include "dff_seq.sv"       // Defines sequence
`include "dff_seqr.sv"      // Defines sequencer
`include "dff_drv.sv"       // Defines driver
`include "dff_mon.sv"       // Defines monitor
`include "dff_scbd.sv"      // Defines scoreboard
`include "dff_agt.sv"       // Defines agent
`include "dff_env.sv"       // Defines environment
`include "dff_test.sv"      // Defines test and runs the environment
